`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:45:33 11/05/2015 
// Design Name: 
// Module Name:    Anti_jitter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Anti_jitter(
    input clk,
    input [3:0] button,
    input [7:0] SW,
    output [3:0] button_out,
    output rst,
    output [3:0] button_pulse,
    output [7:0] SW_OK
    );


endmodule
